module add (
    input a,
    input b,
    output  c
);
assign c = a + b;//666
endmodule